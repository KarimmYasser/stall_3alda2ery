-- Move your existing fetch testbench here
-- (If you have one, copy its contents here)
