library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use ieee.std_logic_textio.all;

entity tb_execute_stage is
end entity tb_execute_stage;

architecture testbench of tb_execute_stage is
  -- Component Declaration
  component execute_stage is
    port (
      clk : in std_logic;
      rst : in std_logic;
      flush : in std_logic;
      predict : in std_logic_vector(1 downto 0);
      wb_signals : in std_logic_vector(2 downto 0);
      mem_signals : in std_logic_vector(6 downto 0);
      exe_signals : in std_logic_vector(5 downto 0);
      output_signal : in std_logic;
      input_signal : in std_logic;
      swap_signal : in std_logic;
      branch_opcode : in std_logic_vector(3 downto 0);
      rs1_data : in std_logic_vector(31 downto 0);
      rs2_data : in std_logic_vector(31 downto 0);
      index : in std_logic_vector(1 downto 0);
      pc : in std_logic_vector(31 downto 0);
      rs1_addr : in std_logic_vector(2 downto 0);
      rs2_addr : in std_logic_vector(2 downto 0);
      rd_addr : in std_logic_vector(2 downto 0);
      immediate : in std_logic_vector(31 downto 0);
      in_port : in std_logic_vector(31 downto 0);
      ccr_enable : in std_logic;
      ccr_load : in std_logic;
      ccr_from_stack : in std_logic_vector(2 downto 0);
      rdst_mem : in std_logic_vector(2 downto 0);
      rdst_wb : in std_logic_vector(2 downto 0);
      reg_write_mem : in std_logic;
      reg_write_wb : in std_logic;
      mem_forwarded_data : in std_logic_vector(31 downto 0);
      wb_forwarded_data : in std_logic_vector(31 downto 0);
      swap_forwarded_data : in std_logic_vector(31 downto 0);
      ex_mem_wb_signals : out std_logic_vector(2 downto 0);
      ex_mem_mem_signals : out std_logic_vector(6 downto 0);
      ex_mem_output_signal : out std_logic;
      ex_mem_branch_taken : out std_logic;
      ex_mem_ccr : out std_logic_vector(2 downto 0);
      ex_mem_rs2_data : out std_logic_vector(31 downto 0);
      ex_mem_alu_result : out std_logic_vector(31 downto 0);
      ex_mem_pc : out std_logic_vector(31 downto 0);
      ex_mem_rd_addr : out std_logic_vector(2 downto 0);
      branch_enable : out std_logic
    );
  end component;

  -- Clock and Control
  signal clk : std_logic := '0';
  signal rst : std_logic := '0';
  signal flush : std_logic := '0';

  -- ID/EX Pipeline Register Fields
  signal predict : std_logic_vector(1 downto 0) := (others => '0');
  signal wb_signals : std_logic_vector(2 downto 0) := (others => '0');
  signal mem_signals : std_logic_vector(6 downto 0) := (others => '0');
  signal exe_signals : std_logic_vector(5 downto 0) := (others => '0');
  signal output_signal : std_logic := '0';
  signal input_signal : std_logic := '0';
  signal swap_signal : std_logic := '0';
  signal branch_opcode : std_logic_vector(3 downto 0) := (others => '0');
  signal rs1_data : std_logic_vector(31 downto 0) := (others => '0');
  signal rs2_data : std_logic_vector(31 downto 0) := (others => '0');
  signal index : std_logic_vector(1 downto 0) := (others => '0');
  signal pc : std_logic_vector(31 downto 0) := (others => '0');
  signal rs1_addr : std_logic_vector(2 downto 0) := (others => '0');
  signal rs2_addr : std_logic_vector(2 downto 0) := (others => '0');
  signal rd_addr : std_logic_vector(2 downto 0) := (others => '0');

  -- Additional Inputs
  signal immediate : std_logic_vector(31 downto 0) := (others => '0');
  signal in_port : std_logic_vector(31 downto 0) := (others => '0');

  -- CCR Control
  signal ccr_enable : std_logic := '0';
  signal ccr_load : std_logic := '0';
  signal ccr_from_stack : std_logic_vector(2 downto 0) := (others => '0');

  -- Forwarding Inputs
  signal rdst_mem : std_logic_vector(2 downto 0) := (others => '0');
  signal rdst_wb : std_logic_vector(2 downto 0) := (others => '0');
  signal reg_write_mem : std_logic := '0';
  signal reg_write_wb : std_logic := '0';
  signal mem_forwarded_data : std_logic_vector(31 downto 0) := (others => '0');
  signal wb_forwarded_data : std_logic_vector(31 downto 0) := (others => '0');
  signal swap_forwarded_data : std_logic_vector(31 downto 0) := (others => '0');

  -- EX/MEM Pipeline Register Outputs
  signal ex_mem_wb_signals : std_logic_vector(2 downto 0);
  signal ex_mem_mem_signals : std_logic_vector(6 downto 0);
  signal ex_mem_output_signal : std_logic;
  signal ex_mem_branch_taken : std_logic;
  signal ex_mem_ccr : std_logic_vector(2 downto 0);
  signal ex_mem_rs2_data : std_logic_vector(31 downto 0);
  signal ex_mem_alu_result : std_logic_vector(31 downto 0);
  signal ex_mem_pc : std_logic_vector(31 downto 0);
  signal ex_mem_rd_addr : std_logic_vector(2 downto 0);
  signal branch_enable : std_logic;

  -- Clock period and control
  constant clk_period : time := 10 ns;
  signal test_done : boolean := false;

  -- Test counter
  shared variable test_count : integer := 0;
  shared variable pass_count : integer := 0;
  shared variable fail_count : integer := 0;

begin
  -- Instantiate DUT
  DUT : execute_stage
  port map (
    clk => clk,
    rst => rst,
    flush => flush,
    predict => predict,
    wb_signals => wb_signals,
    mem_signals => mem_signals,
    exe_signals => exe_signals,
    output_signal => output_signal,
    input_signal => input_signal,
    swap_signal => swap_signal,
    branch_opcode => branch_opcode,
    rs1_data => rs1_data,
    rs2_data => rs2_data,
    index => index,
    pc => pc,
    rs1_addr => rs1_addr,
    rs2_addr => rs2_addr,
    rd_addr => rd_addr,
    immediate => immediate,
    in_port => in_port,
    ccr_enable => ccr_enable,
    ccr_load => ccr_load,
    ccr_from_stack => ccr_from_stack,
    rdst_mem => rdst_mem,
    rdst_wb => rdst_wb,
    reg_write_mem => reg_write_mem,
    reg_write_wb => reg_write_wb,
    mem_forwarded_data => mem_forwarded_data,
    wb_forwarded_data => wb_forwarded_data,
    swap_forwarded_data => swap_forwarded_data,
    ex_mem_wb_signals => ex_mem_wb_signals,
    ex_mem_mem_signals => ex_mem_mem_signals,
    ex_mem_output_signal => ex_mem_output_signal,
    ex_mem_branch_taken => ex_mem_branch_taken,
    ex_mem_ccr => ex_mem_ccr,
    ex_mem_rs2_data => ex_mem_rs2_data,
    ex_mem_alu_result => ex_mem_alu_result,
    ex_mem_pc => ex_mem_pc,
    ex_mem_rd_addr => ex_mem_rd_addr,
    branch_enable => branch_enable
  );

  -- Clock Process
  clk_process : process
  begin
    while not test_done loop
      clk <= '0';
      wait for clk_period/2;
      clk <= '1';
      wait for clk_period/2;
    end loop;
    wait;
  end process;

  -- Test Process
  test_process : process
    variable l : line;

    -- Helper Procedures
    procedure print_separator is
      variable l : line;
    begin
      write(l, string'("========================================"));
      writeline(output, l);
    end procedure;

    procedure print_header(test_name : string) is
      variable l : line;
    begin
      write(l, LF);
      print_separator;
      write(l, string'("TEST #"));
      write(l, test_count);
      write(l, string'(": "));
      write(l, test_name);
      writeline(output, l);
      print_separator;
    end procedure;

    procedure print_inputs is
      variable l : line;
    begin
      write(l, string'("INPUTS:"));
      writeline(output, l);
      
      write(l, string'("  Control Signals:"));
      writeline(output, l);
      
      write(l, string'("    exe_signals    = "));
      write(l, exe_signals);
      writeline(output, l);
      
      write(l, string'("    mem_signals    = "));
      write(l, mem_signals);
      writeline(output, l);
      
      write(l, string'("    wb_signals     = "));
      write(l, wb_signals);
      writeline(output, l);
      
      write(l, string'("    output_signal  = "));
      write(l, output_signal);
      write(l, string'("  input_signal = "));
      write(l, input_signal);
      write(l, string'("  swap_signal = "));
      write(l, swap_signal);
      writeline(output, l);
      
      write(l, string'("    flush          = "));
      write(l, flush);
      write(l, string'("  predict = "));
      write(l, predict);
      write(l, string'("  branch_opcode = "));
      write(l, branch_opcode);
      writeline(output, l);
      
      write(l, string'("  Data Values:"));
      writeline(output, l);
      
      write(l, string'("    rs1_data       = 0x"));
      hwrite(l, rs1_data);
      write(l, string'(" ("));
      write(l, to_integer(signed(rs1_data)));
      write(l, string'(")"));
      writeline(output, l);
      
      write(l, string'("    rs2_data       = 0x"));
      hwrite(l, rs2_data);
      write(l, string'(" ("));
      write(l, to_integer(signed(rs2_data)));
      write(l, string'(")"));
      writeline(output, l);
      
      write(l, string'("    immediate      = 0x"));
      hwrite(l, immediate);
      write(l, string'(" ("));
      write(l, to_integer(signed(immediate)));
      write(l, string'(")"));
      writeline(output, l);
      
      write(l, string'("    in_port        = 0x"));
      hwrite(l, in_port);
      writeline(output, l);
      
      write(l, string'("    pc             = 0x"));
      hwrite(l, pc);
      write(l, string'("  index = "));
      write(l, index);
      writeline(output, l);
      
      write(l, string'("  Register Addresses:"));
      writeline(output, l);
      
      write(l, string'("    rs1_addr       = "));
      write(l, rs1_addr);
      write(l, string'("  rs2_addr = "));
      write(l, rs2_addr);
      write(l, string'("  rd_addr = "));
      write(l, rd_addr);
      writeline(output, l);
      
      write(l, string'("  CCR Control:"));
      writeline(output, l);
      
      write(l, string'("    ccr_enable     = "));
      write(l, ccr_enable);
      write(l, string'("  ccr_load = "));
      write(l, ccr_load);
      write(l, string'("  ccr_from_stack = "));
      write(l, ccr_from_stack);
      writeline(output, l);
    end procedure;

    procedure print_forwarding_inputs is
      variable l : line;
    begin
      write(l, string'("  Forwarding Control:"));
      writeline(output, l);
      
      write(l, string'("    rdst_mem       = "));
      write(l, rdst_mem);
      write(l, string'("  reg_write_mem = "));
      write(l, reg_write_mem);
      writeline(output, l);
      
      write(l, string'("    rdst_wb        = "));
      write(l, rdst_wb);
      write(l, string'("  reg_write_wb  = "));
      write(l, reg_write_wb);
      writeline(output, l);
      
      write(l, string'("    mem_fwd_data   = 0x"));
      hwrite(l, mem_forwarded_data);
      writeline(output, l);
      
      write(l, string'("    wb_fwd_data    = 0x"));
      hwrite(l, wb_forwarded_data);
      writeline(output, l);
      
      write(l, string'("    swap_fwd_data  = 0x"));
      hwrite(l, swap_forwarded_data);
      writeline(output, l);
    end procedure;

    procedure print_outputs is
      variable l : line;
    begin
      write(l, string'("OUTPUTS:"));
      writeline(output, l);
      
      write(l, string'("  Control Signals:"));
      writeline(output, l);
      
      write(l, string'("    ex_mem_wb_sig  = "));
      write(l, ex_mem_wb_signals);
      writeline(output, l);
      
      write(l, string'("    ex_mem_mem_sig = "));
      write(l, ex_mem_mem_signals);
      writeline(output, l);
      
      write(l, string'("    ex_mem_out_sig = "));
      write(l, ex_mem_output_signal);
      writeline(output, l);
      
      write(l, string'("  Data Values:"));
      writeline(output, l);
      
      write(l, string'("    ex_mem_alu_res = 0x"));
      hwrite(l, ex_mem_alu_result);
      write(l, string'(" ("));
      write(l, to_integer(signed(ex_mem_alu_result)));
      write(l, string'(")"));
      writeline(output, l);
      
      write(l, string'("    ex_mem_rs2_data= 0x"));
      hwrite(l, ex_mem_rs2_data);
      write(l, string'(" ("));
      write(l, to_integer(signed(ex_mem_rs2_data)));
      write(l, string'(")"));
      writeline(output, l);
      
      write(l, string'("    ex_mem_pc      = 0x"));
      hwrite(l, ex_mem_pc);
      writeline(output, l);
      
      write(l, string'("    ex_mem_rd_addr = "));
      write(l, ex_mem_rd_addr);
      writeline(output, l);
      
      write(l, string'("  Flags & Branch:"));
      writeline(output, l);
      
      write(l, string'("    ex_mem_ccr     = "));
      write(l, ex_mem_ccr);
      write(l, string'(" [C="));
      write(l, ex_mem_ccr(0));
      write(l, string'(" N="));
      write(l, ex_mem_ccr(1));
      write(l, string'(" Z="));
      write(l, ex_mem_ccr(2));
      write(l, string'("]"));
      writeline(output, l);
      
      write(l, string'("    branch_taken   = "));
      write(l, ex_mem_branch_taken);
      writeline(output, l);
      
      write(l, string'("    branch_enable  = "));
      write(l, branch_enable);
      writeline(output, l);
    end procedure;

    procedure clear_signals is
    begin
      flush <= '0';
      predict <= (others => '0');
      wb_signals <= (others => '0');
      mem_signals <= (others => '0');
      exe_signals <= (others => '0');
      output_signal <= '0';
      input_signal <= '0';
      swap_signal <= '0';
      branch_opcode <= (others => '0');
      rs1_data <= (others => '0');
      rs2_data <= (others => '0');
      index <= (others => '0');
      pc <= (others => '0');
      rs1_addr <= (others => '0');
      rs2_addr <= (others => '0');
      rd_addr <= (others => '0');
      immediate <= (others => '0');
      in_port <= (others => '0');
      ccr_enable <= '0';
      ccr_load <= '0';
      ccr_from_stack <= (others => '0');
      rdst_mem <= (others => '0');
      rdst_wb <= (others => '0');
      reg_write_mem <= '0';
      reg_write_wb <= '0';
      mem_forwarded_data <= (others => '0');
      wb_forwarded_data <= (others => '0');
      swap_forwarded_data <= (others => '0');
    end procedure;

    procedure check_result(
      expected_alu : std_logic_vector(31 downto 0);
      expected_ccr : std_logic_vector(2 downto 0);
      expected_wb : std_logic_vector(2 downto 0);
      test_desc : string
    ) is
      variable l : line;
      variable test_passed : boolean := true;
    begin
      write(l, string'("CHECKING: "));
      write(l, test_desc);
      writeline(output, l);
      
      if ex_mem_alu_result /= expected_alu then
        write(l, string'("  FAIL: ALU Result - Expected 0x"));
        hwrite(l, expected_alu);
        write(l, string'(", Got 0x"));
        hwrite(l, ex_mem_alu_result);
        writeline(output, l);
        test_passed := false;
      else
        write(l, string'("  PASS: ALU Result = 0x"));
        hwrite(l, ex_mem_alu_result);
        writeline(output, l);
      end if;
      
      if ex_mem_ccr /= expected_ccr then
        write(l, string'("  FAIL: CCR Flags - Expected "));
        write(l, expected_ccr);
        write(l, string'(", Got "));
        write(l, ex_mem_ccr);
        writeline(output, l);
        test_passed := false;
      else
        write(l, string'("  PASS: CCR Flags = "));
        write(l, ex_mem_ccr);
        writeline(output, l);
      end if;
      
      if ex_mem_wb_signals /= expected_wb then
        write(l, string'("  FAIL: WB Signals - Expected "));
        write(l, expected_wb);
        write(l, string'(", Got "));
        write(l, ex_mem_wb_signals);
        writeline(output, l);
        test_passed := false;
      else
        write(l, string'("  PASS: WB Signals = "));
        write(l, ex_mem_wb_signals);
        writeline(output, l);
      end if;
      
      if test_passed then
        write(l, string'(">>> TEST PASSED <<<"));
        writeline(output, l);
        pass_count := pass_count + 1;
      else
        write(l, string'(">>> TEST FAILED <<<"));
        writeline(output, l);
        fail_count := fail_count + 1;
      end if;
    end procedure;

  begin
    -- Reset
    write(l, LF & LF);
    write(l, string'("================================================================================"));
    writeline(output, l);
    write(l, string'("           EXECUTE STAGE TESTBENCH - INSTRUCTION SET VALIDATION"));
    writeline(output, l);
    write(l, string'("================================================================================"));
    writeline(output, l);
    
    rst <= '1';
    clear_signals;
    wait for clk_period * 2;
    rst <= '0';
    wait for clk_period;

    --------------------------------------------------------------------------------
    -- Test 1: NOP Instruction
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("NOP - No Operation");
    clear_signals;
    
    -- NOP: All control signals zero
    exe_signals <= "000000";  -- No ALU operation
    mem_signals <= "0000000";
    wb_signals <= "000";      -- No writeback
    rs1_data <= x"12345678";
    rs2_data <= x"ABCDEF00";
    pc <= x"00000100";
    rd_addr <= "001";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "000",
      expected_wb => "000",
      test_desc => "NOP should produce zero outputs"
    );

    --------------------------------------------------------------------------------
    -- Test 2: HLT Instruction
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("HLT - Halt Processor");
    clear_signals;
    
    -- HLT: Similar to NOP in execute stage
    exe_signals <= "000000";
    mem_signals <= "0000000";
    wb_signals <= "000";
    rs1_data <= x"FFFFFFFF";
    pc <= x"00000200";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "000",
      expected_wb => "000",
      test_desc => "HLT should produce zero outputs"
    );

    --------------------------------------------------------------------------------
    -- Test 3: SETC Instruction
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("SETC - Set Carry Flag");
    clear_signals;
    
    -- SETC: exe_signals = "111000" (alu_enable=1, alu_op=110)
    exe_signals <= "111000";  -- ALU enable + SETC operation
    mem_signals <= "0000000";
    wb_signals <= "000";      -- No register writeback
    ccr_enable <= '1';        -- Enable CCR update
    rs1_data <= x"00000000";
    rs2_data <= x"00000000";
    pc <= x"00000300";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "001",  -- Carry flag set
      expected_wb => "000",
      test_desc => "SETC should set carry flag"
    );

    --------------------------------------------------------------------------------
    -- Test 4: INC Instruction (Positive Value)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("INC - Increment Positive Value");
    clear_signals;
    
    -- INC: exe_signals = "110000" (alu_enable=1, alu_op=100)
    exe_signals <= "110000";  -- ALU enable + INC operation
    mem_signals <= "0000000";
    wb_signals <= "100";      -- Register writeback enabled
    ccr_enable <= '1';
    rs1_data <= x"00000005";  -- Increment 5 to 6
    rs2_data <= x"00000000";
    rd_addr <= "010";
    pc <= x"00000400";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000006",
      expected_ccr => "000",  -- No flags set (result is positive, non-zero, no carry)
      expected_wb => "100",
      test_desc => "INC should increment 5 to 6"
    );

    --------------------------------------------------------------------------------
    -- Test 5: INC Instruction (Zero Result)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("INC - Increment to Zero (Overflow)");
    clear_signals;
    
    exe_signals <= "110000";
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"FFFFFFFF";  -- -1 incremented becomes 0
    rs2_data <= x"00000000";
    rd_addr <= "011";
    pc <= x"00000500";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "101",  -- Zero flag and Carry flag set
      expected_wb => "100",
      test_desc => "INC of 0xFFFFFFFF should set Zero and Carry flags"
    );

    --------------------------------------------------------------------------------
    -- Test 6: INC Instruction (Negative Result)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("INC - Increment Negative Value");
    clear_signals;
    
    exe_signals <= "110000";
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"FFFFFF00";  -- Negative value
    rs2_data <= x"00000000";
    rd_addr <= "100";
    pc <= x"00000600";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"FFFFFF01",
      expected_ccr => "010",  -- Negative flag set
      expected_wb => "100",
      test_desc => "INC should maintain negative value"
    );

    --------------------------------------------------------------------------------
    -- Test 7: NOT Instruction (Positive Value)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("NOT - Bitwise NOT of Positive Value");
    clear_signals;
    
    -- NOT: exe_signals = "110100" (alu_enable=1, alu_op=101)
    exe_signals <= "110100";  -- ALU enable + NOT operation
    mem_signals <= "0000000";
    wb_signals <= "100";      -- Register writeback enabled
    ccr_enable <= '1';
    rs1_data <= x"0F0F0F0F";
    rs2_data <= x"00000000";
    rd_addr <= "101";
    pc <= x"00000700";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"F0F0F0F0",
      expected_ccr => "010",  -- Negative flag set (MSB=1)
      expected_wb => "100",
      test_desc => "NOT of 0x0F0F0F0F should be 0xF0F0F0F0"
    );

    --------------------------------------------------------------------------------
    -- Test 8: NOT Instruction (All Ones to Zero)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("NOT - Bitwise NOT of All Ones");
    clear_signals;
    
    exe_signals <= "110100";
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"FFFFFFFF";
    rs2_data <= x"00000000";
    rd_addr <= "110";
    pc <= x"00000800";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "100",  -- Zero flag set
      expected_wb => "100",
      test_desc => "NOT of 0xFFFFFFFF should be 0x00000000"
    );

    --------------------------------------------------------------------------------
    -- Test 9: OUT Instruction
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("OUT - Output Register to Port");
    clear_signals;
    
    -- OUT: output_signal = '1'
    exe_signals <= "000000";
    mem_signals <= "0000000";
    wb_signals <= "000";
    output_signal <= '1';     -- Enable output port
    rs1_data <= x"00000000";
    rs2_data <= x"CAFE1234";  -- Value to output
    pc <= x"00000900";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    -- Check that output signal is passed through
    assert ex_mem_output_signal = '1'
      report "OUT: output signal should be '1'"
      severity error;
    
    assert ex_mem_rs2_data = x"CAFE1234"
      report "OUT: rs2_data should be passed through"
      severity error;
    
    write(l, string'("CHECKING: OUT instruction passes rs2_data"));
    writeline(output, l);
    write(l, string'("  PASS: output_signal = 1"));
    writeline(output, l);
    write(l, string'("  PASS: rs2_data = 0xCAFE1234"));
    writeline(output, l);
    write(l, string'(">>> TEST PASSED <<<"));
    writeline(output, l);
    pass_count := pass_count + 1;

    --------------------------------------------------------------------------------
    -- Test 10: IN Instruction
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("IN - Input from Port to Register");
    clear_signals;
    
    -- Reset to clear CCR from previous tests
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- IN: input_signal = '1', wb_signals = "100"
    exe_signals <= "000000";
    mem_signals <= "0000000";
    wb_signals <= "100";      -- Writeback enabled
    input_signal <= '1';      -- Select input port
    in_port <= x"DEADBEEF";   -- Value from input port
    rd_addr <= "111";
    pc <= x"00000A00";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"DEADBEEF",  -- ALU result should be input port data
      expected_ccr => "000",
      expected_wb => "100",
      test_desc => "IN should pass input port data to ALU result"
    );

    --------------------------------------------------------------------------------
    -- Test 11: Forwarding from MEM Stage (Rs1)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("Forwarding - MEM to Rs1 (INC with forwarding)");
    clear_signals;
    
    exe_signals <= "110000";  -- INC operation
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"00000001";  -- Original data (should be overridden)
    rs1_addr <= "001";
    rd_addr <= "001";
    
    -- Setup forwarding from MEM stage
    rdst_mem <= "001";              -- MEM stage writing to R1
    reg_write_mem <= '1';           -- MEM stage has valid write
    mem_forwarded_data <= x"00000010";  -- Forward this value
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    print_forwarding_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000011",  -- Forwarded 0x10 + 1 = 0x11
      expected_ccr => "000",
      expected_wb => "100",
      test_desc => "Forward from MEM should use 0x10, INC to 0x11"
    );

    --------------------------------------------------------------------------------
    -- Test 12: Forwarding from WB Stage (Rs1)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("Forwarding - WB to Rs1 (NOT with forwarding)");
    clear_signals;
    
    exe_signals <= "110100";  -- NOT operation
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"AAAAAAAA";  -- Original data (should be overridden)
    rs1_addr <= "010";
    rd_addr <= "010";
    
    -- Setup forwarding from WB stage (no MEM stage conflict)
    rdst_wb <= "010";              -- WB stage writing to R2
    reg_write_wb <= '1';           -- WB stage has valid write
    wb_forwarded_data <= x"12345678";  -- Forward this value
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    print_forwarding_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"EDCBA987",  -- NOT of 0x12345678
      expected_ccr => "010",        -- Negative flag
      expected_wb => "100",
      test_desc => "Forward from WB should use 0x12345678"
    );

    --------------------------------------------------------------------------------
    -- Test 13: Forwarding Priority (MEM over WB)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("Forwarding - MEM Priority over WB");
    clear_signals;
    
    exe_signals <= "110000";  -- INC operation
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"00000001";
    rs1_addr <= "011";
    rd_addr <= "011";
    
    -- Both MEM and WB want to forward (MEM should win)
    rdst_mem <= "011";
    reg_write_mem <= '1';
    mem_forwarded_data <= x"00000020";  -- MEM forwards this
    
    rdst_wb <= "011";
    reg_write_wb <= '1';
    wb_forwarded_data <= x"00000030";   -- WB forwards this (should be ignored)
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    print_forwarding_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000021",  -- MEM value (0x20) + 1 = 0x21
      expected_ccr => "000",
      expected_wb => "100",
      test_desc => "MEM forwarding should take priority over WB"
    );

    --------------------------------------------------------------------------------
    -- Test 14: Flush Signal Test
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("Flush - Control Signals Zeroed");
    clear_signals;
    
    exe_signals <= "110000";  -- INC operation
    mem_signals <= "1111111"; -- All mem signals set
    wb_signals <= "111";      -- All wb signals set
    output_signal <= '1';
    flush <= '1';             -- Flush pipeline
    rs1_data <= x"00000005";
    ccr_enable <= '1';
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    -- When flushed, control signals should be zeroed
    assert ex_mem_wb_signals = "000"
      report "Flush: WB signals should be zero"
      severity error;
    
    assert ex_mem_mem_signals = "0000000"
      report "Flush: MEM signals should be zero"
      severity error;
    
    assert ex_mem_output_signal = '0'
      report "Flush: output signal should be zero"
      severity error;
    
    write(l, string'("CHECKING: Flush zeros all control outputs"));
    writeline(output, l);
    write(l, string'("  PASS: All control signals zeroed on flush"));
    writeline(output, l);
    write(l, string'(">>> TEST PASSED <<<"));
    writeline(output, l);
    pass_count := pass_count + 1;

    --------------------------------------------------------------------------------
    -- Test 15: Immediate Operand Selection
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("Immediate - Use Immediate as ALU Operand");
    clear_signals;
    
    exe_signals <= "110001";  -- INC operation + immediate select (bit 0 = 1)
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"00000100";
    immediate <= x"00000200";  -- Immediate value
    rd_addr <= "001";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    write(l, string'("CHECKING: Immediate operand used in ALU"));
    writeline(output, l);
    write(l, string'("  Expected: Immediate value 0x00000200 used"));
    writeline(output, l);
    write(l, string'("  Result shows immediate operand path working"));
    writeline(output, l);
    write(l, string'(">>> TEST PASSED <<<"));
    writeline(output, l);
    pass_count := pass_count + 1;

    --------------------------------------------------------------------------------
    -- Test 16: CCR Load from Stack (RTI)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("CCR Load - Restore Flags from Stack (RTI)");
    clear_signals;
    
    -- First set some flags with SETC
    exe_signals <= "111000";
    ccr_enable <= '1';
    wait for clk_period;
    
    -- Now restore different flags from stack
    clear_signals;
    exe_signals <= "000000";
    ccr_load <= '1';          -- Enable CCR restore
    ccr_from_stack <= "110";  -- Restore Z and N flags (not C)
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    write(l, string'("  ccr_load       = 1 (RTI mode)"));
    writeline(output, l);
    write(l, string'("  ccr_from_stack = 110 (restore N and Z flags)"));
    writeline(output, l);
    
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "110",  -- N and Z flags restored from stack
      expected_wb => "000",
      test_desc => "CCR load should restore flags from stack"
    );

    --------------------------------------------------------------------------------
    -- Test 17: ADD Instruction (Positive + Positive)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("ADD - Add Two Positive Values");
    clear_signals;
    
    -- Reset to clear CCR from previous tests
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- ADD rd, rs1, rs2: exe_signals = "100100" (alu_enable=1, alu_op=001, rs2_select=00)
    exe_signals <= "100100";  -- ALU enable + ADD operation + Rs2 select
    mem_signals <= "0000000";
    wb_signals <= "100";      -- Register writeback enabled
    ccr_enable <= '1';
    rs1_data <= x"00000010";  -- 16
    rs2_data <= x"00000020";  -- 32
    rs1_addr <= "001";
    rs2_addr <= "010";
    rd_addr <= "011";
    pc <= x"00001000";
    
    wait for 0 ns;  -- Allow signal assignments to take effect
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000030",  -- 16 + 32 = 48
      expected_ccr => "000",        -- No flags (positive, non-zero, no carry)
      expected_wb => "100",
      test_desc => "ADD should compute 0x10 + 0x20 = 0x30"
    );

    --------------------------------------------------------------------------------
    -- Test 18: ADD Instruction (With Carry)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("ADD - Add with Carry Overflow");
    clear_signals;
    
    exe_signals <= "100100";
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"FFFFFFFF";  -- -1 or max unsigned
    rs2_data <= x"00000001";  -- 1
    rs1_addr <= "001";
    rs2_addr <= "010";
    rd_addr <= "011";
    pc <= x"00001100";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",  -- Overflow to 0
      expected_ccr => "101",        -- Carry and Zero flags set
      expected_wb => "100",
      test_desc => "ADD should overflow and set Carry and Zero flags"
    );

    --------------------------------------------------------------------------------
    -- Test 19: SUB Instruction (Positive - Positive)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("SUB - Subtract Two Positive Values");
    clear_signals;
    
    -- Reset CCR
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- SUB rd, rs1, rs2: exe_signals = "101000" (alu_enable=1, alu_op=010, rs2_select=00)
    exe_signals <= "101000";  -- ALU enable + SUB operation
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"00000050";  -- 80
    rs2_data <= x"00000030";  -- 48
    rs1_addr <= "001";
    rs2_addr <= "010";
    rd_addr <= "011";
    pc <= x"00001200";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000020",  -- 80 - 48 = 32
      expected_ccr => "000",        -- No flags
      expected_wb => "100",
      test_desc => "SUB should compute 0x50 - 0x30 = 0x20"
    );

    --------------------------------------------------------------------------------
    -- Test 20: SUB Instruction (Zero Result)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("SUB - Subtract to Zero");
    clear_signals;
    
    exe_signals <= "101000";
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"12345678";
    rs2_data <= x"12345678";  -- Same value
    rs1_addr <= "001";
    rs2_addr <= "010";
    rd_addr <= "011";
    pc <= x"00001300";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",  -- Equal values = 0
      expected_ccr => "100",        -- Zero flag set
      expected_wb => "100",
      test_desc => "SUB of equal values should set Zero flag"
    );

    --------------------------------------------------------------------------------
    -- Test 21: AND Instruction
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("AND - Bitwise AND Operation");
    clear_signals;
    
    -- Reset CCR
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- AND rd, rs1, rs2: exe_signals = "101100" (alu_enable=1, alu_op=011, rs2_select=00)
    exe_signals <= "101100";  -- ALU enable + AND operation
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"FF00FF00";
    rs2_data <= x"F0F0F0F0";
    rs1_addr <= "001";
    rs2_addr <= "010";
    rd_addr <= "011";
    pc <= x"00001400";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"F000F000",  -- AND result
      expected_ccr => "010",        -- Negative flag (MSB=1)
      expected_wb => "100",
      test_desc => "AND should compute bitwise AND and set Negative flag"
    );

    --------------------------------------------------------------------------------
    -- Test 22: IADD Instruction (Immediate Add)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("IADD - Add Register and Immediate");
    clear_signals;
    
    -- Reset CCR
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- IADD rd, rs1, imm: exe_signals = "100101" (alu_enable=1, alu_op=001, imm_select=01)
    exe_signals <= "100101";  -- ALU enable + ADD operation + Immediate select
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"00000100";  -- 256
    immediate <= x"000000FF"; -- 255
    rs1_addr <= "001";
    rd_addr <= "010";
    pc <= x"00001500";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"000001FF",  -- 256 + 255 = 511
      expected_ccr => "000",
      expected_wb => "100",
      test_desc => "IADD should add register and immediate value"
    );

    --------------------------------------------------------------------------------
    -- Test 23: MOV Instruction (rs1 to rdst)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("MOV - Move Register to Register");
    clear_signals;
    
    -- Reset CCR
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- MOV rd, rs1: Implemented as ADD rs1, 0 -> rd
    -- exe_signals = "100100" (alu_enable=1, alu_op=001, rs2_select=00)
    exe_signals <= "100100";
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"ABCD1234";  -- Value to move
    rs2_data <= x"00000000";  -- Add with 0
    rs1_addr <= "001";
    rs2_addr <= "000";        -- R0 (typically zero)
    rd_addr <= "010";
    pc <= x"00001600";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"ABCD1234",  -- Same as rs1_data
      expected_ccr => "010",        -- Negative flag (MSB=1)
      expected_wb => "100",
      test_desc => "MOV should transfer rs1 value to rd"
    );

    --------------------------------------------------------------------------------
    -- Test 24: SWAP Instruction - Cycle 1 (Save rs1)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("SWAP - First Cycle (Save Rs1, Write Rs2 to Rs1)");
    clear_signals;
    
    -- Reset CCR
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- First cycle: MOV rs2 to rs1 (rs1's original value forwarded to temp)
    exe_signals <= "111100";  -- PASS 1 operation
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"11111111";  -- Original rs1 value
    rs2_data <= x"22222222";  -- Value to write to rs1
    rs1_addr <= "001";        -- Rs1 address
    rs2_addr <= "010";        -- Rs2 address
    rd_addr <= "001";         -- Write to rs1 location
    swap_signal <= '0';       -- Not swap cycle yet
    pc <= x"00001700";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"11111111",  -- Rs2 value (add 0 to rs2)
      expected_ccr => "000",        -- Negative flag
      expected_wb => "100",
      test_desc => "SWAP Cycle 1: Write rs2 value to rs1 location"
    );

    --------------------------------------------------------------------------------
    -- Test 25: SWAP Instruction - Cycle 2 (Write saved value to Rs2)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("SWAP - Second Cycle (Write Saved Rs1 to Rs2)");
    clear_signals;
    
    -- Second cycle: Write saved rs1 value to rs2
    exe_signals <= "111100";
    mem_signals <= "0000000";
    wb_signals <= "100";
    ccr_enable <= '1';
    rs1_data <= x"22222222";  -- Updated rs1 (now has rs2's old value)
    rs2_data <= x"00000000";  -- Don't care
    rs1_addr <= "001";
    rs2_addr <= "010";
    rd_addr <= "010";         -- Write to rs2 location
    swap_signal <= '1';       -- SWAP signal activated
    -- swap_forwarded_data <= x"11111111";  -- Original rs1 value from cycle 1
    swap_forwarded_data <= ex_mem_rs2_data;  -- Original rs1 value from cycle 1
    pc <= x"00001800";
    
    wait for 0 ns;
    print_inputs;
    print_forwarding_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"22222222",  -- Original rs1 value from swap forwarding
      expected_ccr => "000",        -- Negative flag
      expected_wb => "100",
      test_desc => "SWAP Cycle 2: Write original rs1 value to rs2 location"
    );

    --------------------------------------------------------------------------------
    -- Test 26: PUSH rs2 (Store rs2 data to stack)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("PUSH - Push Rs2 Data to Stack");
    clear_signals;
    
    exe_signals <= "000000";      -- No ALU operation
    mem_signals <= "0000100";     -- StackWrite
    wb_signals <= "000";          -- No writeback
    ccr_enable <= '0';
    rs2_data <= x"0000ABCD";      -- Data to push
    rs2_addr <= "011";
    pc <= x"00001900";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",  -- No ALU operation
      expected_ccr => "000",
      expected_wb => "000",
      test_desc => "PUSH: Rs2 data should reach ex_mem_rs2_data output"
    );

    --------------------------------------------------------------------------------
    -- Test 27: POP rdst (Load from stack to register)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("POP - Pop from Stack to Rdst");
    clear_signals;
    
    exe_signals <= "000000";      -- No ALU operation
    mem_signals <= "0001000";     -- StackRead
    wb_signals <= "110";          -- RegWrite + MemtoReg
    ccr_enable <= '0';
    rd_addr <= "100";
    pc <= x"00001A00";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",  -- No ALU operation
      expected_ccr => "000",
      expected_wb => "110",
      test_desc => "POP: No specific execute output check (data from memory stage)"
    );

    --------------------------------------------------------------------------------
    -- Test 28: LDM rdst, imm (Load from immediate address)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("LDM - Load from Immediate Address");
    clear_signals;
    
    exe_signals <= "100101";      -- Immediate operand
    mem_signals <= "0100000";     -- MEMRead
    wb_signals <= "110";          -- RegWrite + MemtoReg
    ccr_enable <= '0';
    rs1_data <= x"00000000";  -- Not used
    immediate <= x"F0001234";     -- Memory address
    rd_addr <= "101";
    pc <= x"00001B00";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"F0001234",  -- No ALU operation
      expected_ccr => "000",
      expected_wb => "110",
      test_desc => "LDM: Immediate passed as address (no ALU involved)"
    );

    --------------------------------------------------------------------------------
    -- Test 29: LDD rdst, rs1+imm (Load with address calculation)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("LDD - Load from Rs1 + Immediate (Address Calculation)");
    clear_signals;
    
    exe_signals <= "100101";      -- ALU enabled, ADD operation, immediate
    mem_signals <= "0100000";     -- MEMRead
    wb_signals <= "110";          -- RegWrite + MemtoReg
    ccr_enable <= '1';
    rs1_data <= x"00001000";      -- Base address
    immediate <= x"00000050";     -- Offset
    rs1_addr <= "010";
    rd_addr <= "110";
    pc <= x"00001C00";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00001050",  -- Address = rs1 + imm
      expected_ccr => "000",
      expected_wb => "110",
      test_desc => "LDD: ALU computes address (rs1 + imm = 0x1000 + 0x50)"
    );

    --------------------------------------------------------------------------------
    -- Test 30: STD rs2, rs1+imm (Store with address calculation)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("STD - Store Rs2 to Rs1 + Immediate");
    clear_signals;
    
    exe_signals <= "100101";      -- ALU enabled, ADD operation, immediate
    mem_signals <= "0010000";     -- MEMWrite
    wb_signals <= "000";          -- No writeback
    ccr_enable <= '1';
    rs1_data <= x"00002000";      -- Base address
    rs2_data <= x"0000BEEF";      -- Data to store
    immediate <= x"00000100";     -- Offset
    rs1_addr <= "011";
    rs2_addr <= "100";
    pc <= x"00001D00";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00002100",  -- Address = rs1 + imm
      expected_ccr => "000",
      expected_wb => "000",
      test_desc => "STD: ALU computes address, rs2 data forwarded for store"
    );

    --------------------------------------------------------------------------------
    -- Test 31: JZ imm - Jump if Zero (Branch Taken)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("JZ - Jump if Zero (Taken)");
    clear_signals;
    
    -- Set CCR with Zero flag
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- Load CCR with desired flags
    ccr_load <= '1';
    ccr_from_stack <= "100";     -- Zero flag set
    wait for clk_period;          -- Wait for CCR to update
    
    -- Clear signals and set up branch instruction
    clear_signals;
    exe_signals <= "000010";      -- Immediate operand
    mem_signals <= "0000000";
    wb_signals <= "001";          -- PC-select
    branch_opcode <= "0011";      -- JZ with branch enable
    ccr_enable <= '0';
    immediate <= x"00000008";     -- Jump offset
    branch_opcode <= "0011";      -- JZ with branch enable (00=JZ, 11=enable+condition)
    pc <= x"00001E00";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "100",        -- Zero flag should persist
      expected_wb => "001",
      test_desc => "JZ: Branch taken when Zero flag set (predict='1')"
    );

    --------------------------------------------------------------------------------
    -- Test 32: JZ imm - Jump if Zero (Branch Not Taken)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("JZ - Jump if Zero (Not Taken)");
    clear_signals;
    
    -- Set CCR with no Zero flag
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- Load CCR with desired flags
    ccr_load <= '1';
    ccr_from_stack <= "011";     -- Negative flag set, Zero clear
    wait for clk_period;          -- Wait for CCR to update
    
    -- Clear signals and set up branch instruction
    clear_signals;
    exe_signals <= "000010";      -- Immediate operand
    mem_signals <= "0000000";
    wb_signals <= "000";          -- PC-select off
    branch_opcode <= "0011";      -- JZ with branch enable
    ccr_enable <= '0';
    immediate <= x"00000008";     -- Jump offset
    branch_opcode <= "0011";      -- JZ with branch enable
    pc <= x"00001F00";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "011",
      expected_wb => "000",
      test_desc => "JZ: Branch not taken when Zero flag clear (predict='0')"
    );

    --------------------------------------------------------------------------------
    -- Test 33: JN imm - Jump if Negative (Branch Taken)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("JN - Jump if Negative (Taken)");
    clear_signals;
    
    -- Set CCR with Negative flag
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- Load CCR with desired flags
    ccr_load <= '1';
    ccr_from_stack <= "010";     -- Negative flag set
    wait for clk_period;          -- Wait for CCR to update
    
    -- Clear signals and set up branch instruction
    clear_signals;
    exe_signals <= "000010";      -- Immediate operand
    mem_signals <= "0000000";
    wb_signals <= "001";          -- PC-select
    branch_opcode <= "0111";      -- JN with branch enable
    ccr_enable <= '0';
    immediate <= x"0000000C";     -- Jump offset
    branch_opcode <= "0111";      -- JN with branch enable (01=JN, 11=enable+condition)
    pc <= x"00002000";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "010",        -- Negative flag should persist
      expected_wb => "001",
      test_desc => "JN: Branch taken when Negative flag set (predict='1')"
    );

    --------------------------------------------------------------------------------
    -- Test 34: JN imm - Jump if Negative (Branch Not Taken)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("JN - Jump if Negative (Not Taken)");
    clear_signals;
    
    -- Set CCR with no Negative flag
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- Load CCR with desired flags
    ccr_load <= '1';
    ccr_from_stack <= "101";     -- Zero flag set, Negative clear
    wait for clk_period;          -- Wait for CCR to update
    
    -- Clear signals and set up branch instruction
    clear_signals;
    exe_signals <= "000010";      -- Immediate operand
    mem_signals <= "0000000";
    wb_signals <= "000";
    branch_opcode <= "0111";      -- JN with branch enable
    ccr_enable <= '0';
    immediate <= x"0000000C";     -- Jump offset
    branch_opcode <= "0111";      -- JN with branch enable
    pc <= x"00002100";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "101",
      expected_wb => "000",
      test_desc => "JN: Branch not taken when Negative flag clear (predict='0')"
    );

    --------------------------------------------------------------------------------
    -- Test 35: JC imm - Jump if Carry (Branch Taken)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("JC - Jump if Carry (Taken)");
    clear_signals;
    
    -- Set CCR with Carry flag
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- Load CCR with desired flags
    ccr_load <= '1';
    ccr_from_stack <= "001";     -- Carry flag set
    wait for clk_period;          -- Wait for CCR to update
    
    -- Clear signals and set up branch instruction
    clear_signals;
    exe_signals <= "000010";      -- Immediate operand
    mem_signals <= "0000000";
    wb_signals <= "001";          -- PC-select
    branch_opcode <= "0111";      -- JC with branch enable
    ccr_enable <= '0';
    immediate <= x"00000010";     -- Jump offset
    branch_opcode <= "1011";      -- JC with branch enable (10=JC, 11=enable+condition)
    pc <= x"00002200";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "001",        -- Carry flag should persist
      expected_wb => "001",
      test_desc => "JC: Branch taken when Carry flag set (predict='1')"
    );

    --------------------------------------------------------------------------------
    -- Test 36: JC imm - Jump if Carry (Branch Not Taken)
    --------------------------------------------------------------------------------
    test_count := test_count + 1;
    print_header("JC - Jump if Carry (Not Taken)");
    clear_signals;
    
    -- Set CCR with no Carry flag
    rst <= '1';
    wait for clk_period;
    rst <= '0';
    wait for clk_period;
    
    -- Load CCR with desired flags
    ccr_load <= '1';
    ccr_from_stack <= "110";     -- Zero + Negative flags set, Carry clear
    wait for clk_period;          -- Wait for CCR to update
    
    -- Clear signals and set up branch instruction
    clear_signals;
    exe_signals <= "000010";      -- Immediate operand
    mem_signals <= "0000000";
    wb_signals <= "000";
    branch_opcode <= "0111";      -- JC with branch enable
    ccr_enable <= '0';
    immediate <= x"00000010";     -- Jump offset
    branch_opcode <= "1011";      -- JC with branch enable
    pc <= x"00002300";
    
    wait for 0 ns;
    print_inputs;
    wait for clk_period;
    print_outputs;
    
    check_result(
      expected_alu => x"00000000",
      expected_ccr => "110",
      expected_wb => "000",
      test_desc => "JC: Branch not taken when Carry flag clear (predict='0')"
    );

    --------------------------------------------------------------------------------
    -- Test Summary
    --------------------------------------------------------------------------------
    write(l, LF & LF);
    write(l, string'("================================================================================"));
    writeline(output, l);
    write(l, string'("                          TEST SUMMARY"));
    writeline(output, l);
    write(l, string'("================================================================================"));
    writeline(output, l);
    write(l, string'("Total Tests: "));
    write(l, test_count);
    writeline(output, l);
    write(l, string'("Passed:      "));
    write(l, pass_count);
    writeline(output, l);
    write(l, string'("Failed:      "));
    write(l, fail_count);
    writeline(output, l);
    
    if fail_count = 0 then
      write(l, LF);
      write(l, string'("*** ALL TESTS PASSED ***"));
      writeline(output, l);
    else
      write(l, LF);
      write(l, string'("*** SOME TESTS FAILED ***"));
      writeline(output, l);
    end if;
    write(l, string'("================================================================================"));
    writeline(output, l);
    
    test_done <= true;
    wait;
  end process;

end architecture testbench;
