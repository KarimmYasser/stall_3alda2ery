-- Placeholder fetch testbench
-- TODO: Implement fetch stage testbench

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fetch_tb is
end entity fetch_tb;

architecture testbench of fetch_tb is
begin
    -- TODO: Add testbench implementation
end architecture testbench;
